//============================================================
// File: XXX_uvm_env_template.sv
// Description: Generic UVM Environment Template
// Author: Mohamed Essam
//============================================================


//============================================================
// PACKAGE: XXX_shared_pkg
//============================================================


//============================================================
// PACKAGE: XXX_config_pkg
//============================================================


//============================================================
// INTERFACE: XXX_if
//============================================================



//============================================================
// PACKAGE: XXX_seq_item_pkg
//============================================================



//============================================================
// PACKAGE: XXX_main_seq_pkg
//============================================================


//============================================================
// PACKAGE: XXX_rst_seq_pkg
//============================================================



//============================================================
// PACKAGE: XXX_sequencer_pkg
//============================================================



//============================================================
// PACKAGE: XXX_driver_pkg
//============================================================



//============================================================
// PACKAGE: XXX_monitor_pkg
//============================================================



//============================================================
// PACKAGE: XXX_agent_pkg
//============================================================



//============================================================
// PACKAGE: XXX_scoreboard_pkg
//============================================================



//============================================================
// PACKAGE: XXX_coverage_pkg
//============================================================



//============================================================
// PACKAGE: XXX_env_pkg
//============================================================



//============================================================
// PACKAGE: XXX_test_pkg
//============================================================


//============================================================
// END OF FILE
//============================================================

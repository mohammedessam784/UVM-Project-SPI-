import SPI_slave_shared_pkg::*;
module SPI_slave_sva(SPI_slave_if.DUT SPI_slaveif);


endmodule